`default_nettype none

module test;
    // Tiny Tapeout testbench template
    initial begin
        $display("Tiny Tapeout test started.");
        $finish;
    end
endmodule
